-------------------------------------------------------------------------------
-- Title         : 
-- Project       : 
-------------------------------------------------------------------------------
-- File          : edit_msg.vhd
-- Author        : Pedro Messias Jose da Cunha Bastos
-- Company       : 
-- Created       : 2015-04-17
-- Last update   : 2015-05-19
-- Target Device : 
-- Standard      : VHDL'93/02
-------------------------------------------------------------------------------
-- Description   : Edit_msg Implementation
-------------------------------------------------------------------------------
-- Copyright (c) 2015 
-------------------------------------------------------------------------------
-- Revisions     :
-- Date        Version  Author  Description
-- 2015-04-17  1.0      Ordep   Created
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity edit_msg is

  port (
    sysclk  : in std_logic;                    -- global clock
    reset_n : in std_logic);                   -- global reset
  data_o : out std_logic_vector (31 downto 0)  --
    );

end entity edit_msg;

architecture edit_msg_rtl of edit_msg is

  type MSG_ST_TYPE is (ST_INIT);
  type msg is natural range 0 to 7 of std_logic_vector(31 downto 0);

  signal state_reg  : MSG_ST_TYPE;
  signal state_next : MSG_ST_TYPE;

begin  -- architecture edit_msg_rtl

  process(reset_n, sysclk)

  begin

    if reset_n = '0' then
      state_reg <= ST_INIT;

    elsif rising_edge(sysclk) then
      state_reg <= state_next;

    end if;

  end process;


  process (state_reg)

  begin

    state_next <= state_reg;

    case state_reg is

      when ST_INIT =>

    end process;



  end architecture edit_msg_rtl;
























































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































