-------------------------------------------------------------------------------
-- Title         : 
-- Project       : 
-------------------------------------------------------------------------------
-- File          : edit_msg.vhd
-- Author        : Pedro Messias Jose da Cunha Bastos
-- Company       : 
-- Created       : 2015-04-17
-- Last update   : 2015-05-19
-- Target Device : 
-- Standard      : VHDL'93/02
-------------------------------------------------------------------------------
-- Description   : Edit_msg Implementation
-------------------------------------------------------------------------------
-- Copyright (c) 2015 
-------------------------------------------------------------------------------
-- Revisions     :
-- Date        Version  Author  Description
-- 2015-04-17  1.0      Ordep   Created
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity edit_msg is

  port (
    sysclk  : in std_logic;             -- global clock
    reset_n : in std_logic);            -- global reset

end entity edit_msg;

type MSG_ST_TYPE is ();
type msg is natural range 0 to 7 of std_logic_vector(31 downto 0);

architecture edit_msg_rtl of edit_msg is

begin  -- architecture edit_msg_rtl



end architecture edit_msg_rtl;
























































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































